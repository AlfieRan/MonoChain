module memory
import os
import json

pub struct Cache_Struct{
	// Since V does not allow for lists to be map keys, all keys must be json encoded then used as a string key
	pub mut:
		loaded bool
		grudges map[string]i8	// maps a node pub key/id to a local grudge -> negative is good, positive is a bad.
}

pub fn (mut Cache Cache_Struct) load_cache(file_path string){
	data = read_file(file_path, Cache, true)
	// no Trust/grudge file, need to generate a new one
}

pub fn (Cache Cache_Struct) save (file_location string){
	raw := json.encode(Cache)

	os.write_file(file_location, raw) or { // try and write data to file
		// if it failed, run the recursion depth checker to ensure there hasn't been too many failed attempts
		eprintln('Failed to save Trust/Grunge file.')
		exit(1)
	}
}