module utils

pub const (
	confirm = ["y", "yes", "true", "confirm", "affirmative", "1"]
	deny = ["n", "no", "false", "deny", "big no no", "0"]
	alphabet_lower = 97
	alphabet_upper = 122
)