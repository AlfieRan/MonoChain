module configuration
// Use DSA algorithm to generate keys here if the user doesn't have any