module cryptography

type Keys_type = Keys
